`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:14:41 11/03/2017 
// Design Name: 
// Module Name:    MemoryController 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MemoryController(
    );


	// still in VGA controller. Needs to be passed back and fort
	wire req;
	wire [7:0] VGAdata;
	wire [13:0] RAMaddress;
	wire [15:0] RAMdata;
	
	//synthesis attribute box_type VGARAM "black_box"
	VGARAM	_VGARAM(.clka(clk),.addra(RAMaddress),.douta(RAMdata), .wea(1'b0), .dina(16'b0));
endmodule
